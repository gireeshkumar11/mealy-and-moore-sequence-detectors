module seq_detector_mealy_tb;

    reg clk;
    reg reset;
    reg in;
    wire out;
    wire [1:0] currentstate, nextstate;

    seq_detector_mealy dut (
        .in(in),
        .clk(clk),
        .reset(reset),
        .out(out),
        .currentstate(currentstate),
        .nextstate(nextstate)
    );

    always #5 clk = ~clk;

    initial begin
      
        clk = 0;
        reset = 1;
        in = 0;

    
        #10 reset = 0;
        
        #10 in = 1; 
        #10 in = 0;
        #10 in = 0;
        #10 in = 1;   // 1001 detected 
        #10 in = 0;
        #10 in = 0;
        #10 in = 1;   // second 1001 detected

        #20 $finish;
    end
    endmodule
